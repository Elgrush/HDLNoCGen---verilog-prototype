`ifndef _queue_parameters_svh_
`define _queue_parameters_svh_

`include "noc.svh"

`define EN 4 // number of queue entries

`endif
