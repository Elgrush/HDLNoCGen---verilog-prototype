`ifndef _router_parameters_svh_
`define _router_parameters_svh_

`include "noc.svh"

`define REN 5 // number of router entries
`define CS 2 // size of single coordinate part
`define RMS 4 // router marker size

`endif
