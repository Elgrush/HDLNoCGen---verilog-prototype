`ifndef _noc_parameters_svh_
`define _noc_parameters_svh_

`define PL 8// length of datapack
`define CS 2 // size of single coordinate part
`define RMS 4 // router marker size
`define RN 16 // number of routers in network
`define X 4 // number of routers in network on X axis
`define Y 4 // number of routers in network on Y axis
`define CLK_PERIOD 2 // clock period time

`endif
